module seg_disp_top(
	input  [5:0] bin,
	output [6:0] bcd_1, bcd_10
);

	// shift-and-add-3 algorithm
	// THIS IS HARD CODED FOR 6-bit binary input, with 2 digit BCD output
	
	
endmodule
