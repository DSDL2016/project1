module sub_top #(
	parameter width = 6
)(
	input	 [width-1:0] a,
	input  [width-1:0] b,
	output [width-1:0] out,
	output				 overflow
);

endmodule
