module div_top #(
	parameter width = 6
)(
	input						  clk,
	input						  sign,
	input		  [width-1:0] dividend, divider,
	output reg [width-1:0] quotient,
	output	  [width-1:0] remainder,
	output					  ready
);

	
endmodule
